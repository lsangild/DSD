----- Libraries -----
LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-----Package----
package easy is
	constant iBits	: integer;
end easy;

package body easy is
	constant iBits : integer := 8;
end package body easy;