library verilog;
use verilog.vl_types.all;
entity full_adder is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        cin             : in     vl_logic;
        sum             : out    vl_logic;
        cout            : out    vl_logic;
        c1              : out    vl_logic;
        c2              : out    vl_logic;
        s1              : out    vl_logic
    );
end full_adder;
