----- Libraries -----
library ieee;
use ieee.std_logic_1164.all;


entity Mee-Moo is
	port(	
	
	);

end Mee-Moo;